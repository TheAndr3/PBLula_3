module fsm_main (
    input wire clk,                      // Clock de 50MHz
    input wire reset,                    // Reset global
    input wire cmd_iniciar,              // Comando do mestre para iniciar enchimento
    input wire sensor_nivel,             // SW1 - Sensor de nível (1 = cheia)
    input wire alarme_rolha,             // Alarme de falta de rolha
	 input wire aprovado,                // SW2 - Aprovar CQ
    input wire reprovado,              // SW3 - Reprovar CQ
	 output wire esteira,						// LEDR[9] - Motor ligado
    output wire valvula_ativa,           // LEDR[8] - Válvula de enchimento
    output wire vedacao_ativa,           // LEDR[7] - Atuador de vedação
    output wire decrementar_rolha,       // Sinal para decrementar contador
    output wire descarte_ativo,          // LEDR[6] - Atuador de descarte
    output wire garrafa_aprovada,        // Sinal para incrementar contador de dúzias
	 output wire posicao_cq
);

    // Estados da FSM
    localparam IDLE = 4'b0000 ;
	 localparam ESTEIRA = 4'b0001 ;
    localparam ENCHENDO = 4'b0010 ;
    localparam CONCLUIDO = 4'b0011 ;
	 localparam VEDANDO =  4'b0100 ;
	 localparam POSICAO_CQ = 4'b0101 ;
	 localparam DESCARTANDO = 4'b0110 ;
	 localparam APROVADO = 4'b0111 ;
	 
	 reg [25:0] tempo_motor;
	 reg [25:0] tempo_ved;
	 reg [25:0] tempo_descarte;
	 reg [25:0] tempo_aprovado;
	 parameter UM_SEGUNDO = 26'd50000000;
	 reg motor;
    
    reg [3:0] estado_atual;
    
    // Lógica de transição de estados (SEQUENCIAL)
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            estado_atual <= IDLE;
				tempo_motor <= 0;
				tempo_ved <= 0;
				motor <= 1'b0;
				tempo_descarte <= 0;
				tempo_aprovado <= 0;
        end else begin
            case (estado_atual)
                IDLE: begin
							tempo_motor <= 0;
							motor <= 1'b0;
                    if (cmd_iniciar) begin
                        estado_atual <= ESTEIRA;
                    end
                end
					 
					 ESTEIRA: begin
							motor <= 1'b1;
							tempo_motor <= tempo_motor + 1;
							tempo_descarte <= 0;
							tempo_ved <= 0;
							tempo_aprovado <= 0;
							
							if (tempo_motor >= UM_SEGUNDO) begin
								motor <= 1'b0;
								tempo_motor <= 0;
								estado_atual <= ENCHENDO;
							end
                end
                
                ENCHENDO: begin
						  	
                    // Transição ocorre quando sensor de nível detecta garrafa cheia
                    if (sensor_nivel && !alarme_rolha) begin
                        estado_atual <= VEDANDO;
                    end
						  else if (alarme_rolha) begin
								estado_atual <= IDLE;
							end
                end
					 
					 VEDANDO: begin
						tempo_ved <= tempo_ved+1;
						if (tempo_ved >= UM_SEGUNDO) begin
							tempo_ved <= 0;
							estado_atual <= POSICAO_CQ;
						end
					 end
					 
					 POSICAO_CQ: begin
						  
                    if (reprovado && !aprovado) begin
                        estado_atual <= DESCARTANDO;
                    end
						  if (aprovado && !reprovado) begin
                        estado_atual <= APROVADO;
                    end
					 end
                
					 DESCARTANDO: begin
							tempo_descarte <= tempo_descarte+1;
							
							if (tempo_descarte >= UM_SEGUNDO) begin
								tempo_descarte <= 0;
								 estado_atual <= ESTEIRA;
							end
                    
                end
                
                APROVADO: begin
                    tempo_aprovado <= tempo_aprovado+1;
						  
                    if (tempo_aprovado >= UM_SEGUNDO) begin
								tempo_aprovado <= 0;
                        estado_atual <= ESTEIRA;
                    end
						  
                end
                
                default: begin
                    estado_atual <= IDLE;
                end
            endcase
        end
    end
    
    // ========================================================================
    // LÓGICA MOORE: Saídas dependem APENAS do ESTADO (ESTRUTURAL - PORTAS)
    // ========================================================================
    // Extração dos bits do estado (2 bits: estado_atual[1:0])
    // Codificação: IDLE=00, ENCHENDO=01, CONCLUIDO=10
    wire state_bit0, state_bit1, state_bit2, state_bit3;
    buf (state_bit0, estado_atual[0]);
    buf (state_bit1, estado_atual[1]);
	 buf (state_bit2, estado_atual[2]);
	 buf (state_bit3, estado_atual[3]);
    
    // Sinais intermediários
    wire not_state_bit0, not_state_bit1, not_state_bit2, not_state_bit3;
    not (not_state_bit0, state_bit0);
    not (not_state_bit1, state_bit1);
	 not (not_state_bit2, state_bit2);
	 not (not_state_bit3, state_bit3);
	 
	 // Ativação do motor
	 buf (esteira, motor);
    
    // valvula_ativa = 1 quando estado_atual == ENCHENDO (01)
    // Ou seja: state_bit1=0 AND state_bit0=1
    and (valvula_ativa, not_state_bit3, not_state_bit2, state_bit1, not_state_bit0);
	 
	 //Vedaçao ativa
	 wire estado_ved;
	 and (estado_ved, not_state_bit3, state_bit2, not_state_bit1, not_state_bit0);
	 buf (vedacao_ativa , estado_ved);
	 buf (decrementar_rolha, estado_ved);
	 
	 // Estado posicao cq (0101)
	 and (posicao_cq, not_state_bit3, state_bit2, not_state_bit1, state_bit0);
    	 
	 // Estado do descarte (0110)
	 and (descarte_ativo, not_state_bit3, state_bit2, state_bit1, not_state_bit0);
	 
	 // Estado aprovado (0111)
	 and (garrafa_aprovada, not_state_bit3, state_bit2, state_bit1, state_bit0);

endmodule